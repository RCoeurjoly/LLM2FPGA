module matmul_bitstream_top(
  input logic clock,
  input logic reset,
  input logic in3_valid,
  input logic out0_ready,
  input logic in0_ld0_addr_ready,
  input logic in1_ld0_addr_ready,
  output logic in2_st0_done_ready,
  input logic in2_st0_ready,
  input logic [31:0] in0_ld0_data,
  input logic in0_ld0_data_valid,
  input logic [31:0] in1_ld0_data,
  input logic in1_ld0_data_valid,
  output logic [31:0] in2_st0,
  output logic in2_st0_valid,
  output logic in2_st0_done_valid,
  output logic out0_valid,
  output logic [3:0] in0_ld0_addr,
  output logic in0_ld0_addr_valid,
  output logic [3:0] in1_ld0_addr,
  output logic in1_ld0_addr_valid,
  output logic in0_ld0_data_ready,
  output logic in1_ld0_data_ready,
  output logic in3_ready
);

  main u_dut(
    .clock(clock),
    .reset(reset),
    .in3_valid(in3_valid),
    .out0_ready(out0_ready),
    .in0_ld0_addr_ready(in0_ld0_addr_ready),
    .in1_ld0_addr_ready(in1_ld0_addr_ready),
    .in2_st0_ready(in2_st0_ready),
    .in2_st0_done_ready(in2_st0_done_ready),
    .in2_st0_done_valid(in2_st0_done_valid),
    .in2_st0(in2_st0),
    .in2_st0_valid(in2_st0_valid),
    .out0_valid(out0_valid),
    .in0_ld0_addr(in0_ld0_addr),
    .in0_ld0_addr_valid(in0_ld0_addr_valid),
    .in1_ld0_addr(in1_ld0_addr),
    .in1_ld0_addr_valid(in1_ld0_addr_valid),
    .in0_ld0_data(in0_ld0_data),
    .in0_ld0_data_valid(in0_ld0_data_valid),
    .in1_ld0_data(in1_ld0_data),
    .in1_ld0_data_valid(in1_ld0_data_valid),
    .in0_ld0_data_ready(in0_ld0_data_ready),
    .in1_ld0_data_ready(in1_ld0_data_ready),
    .in3_ready(in3_ready)
  );
endmodule
